module dual_port_ram
